library verilog;
use verilog.vl_types.all;
entity Question_1_tb is
end Question_1_tb;
